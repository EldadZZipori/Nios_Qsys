module modulator_signal_selector
# (parameter S = 12)
(
	input logic [7:0] signal_selector,
	input logic [3:0] modulation_selector,
	
	input	logic [11:0]	sin_wave,
	input logic [11:0]	cos_wave,
	input logic [11:0]	squ_wave,
	input	logic [11:0]	saw_wave,
	
	input logic [11:0]	sin_bpsk,
	input logic [11:0]	cos_bpsk,
	input logic [11:0]	squ_bpsk,
	input logic [11:0]	saw_bpsk,
	
	input	logic [11:0]	sin_ask,
	input	logic [11:0]	cos_ask,
	input logic [11:0]	squ_ask,
	input logic [11:0]	saw_ask,

	output logic [11:0] selected_modulation,
	output logic [11:0] selected_signal
);

 /*
	always_comb begin
		case (signal_selector)
			0:
			1:
			2:
			3:
			default:
		endcase
	end
	
	always_comb begin
		case (modulation_selector)
			0:
			1:
			2:
			3:
			default:
		endcase
	end*/
endmodule
